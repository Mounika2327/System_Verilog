module add(
  input [2:0]a,b,
  output [3:0] c );
  assign c= a+b;
endmodule
